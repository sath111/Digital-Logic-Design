library verilog;
use verilog.vl_types.all;
entity SHIFTER1V1_vlg_vec_tst is
end SHIFTER1V1_vlg_vec_tst;
