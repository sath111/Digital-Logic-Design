library verilog;
use verilog.vl_types.all;
entity ABSMINMAX_vlg_vec_tst is
end ABSMINMAX_vlg_vec_tst;
