library verilog;
use verilog.vl_types.all;
entity QUEUERAM_vlg_vec_tst is
end QUEUERAM_vlg_vec_tst;
