library verilog;
use verilog.vl_types.all;
entity ABSMINMAXADDSUB_vlg_vec_tst is
end ABSMINMAXADDSUB_vlg_vec_tst;
