library verilog;
use verilog.vl_types.all;
entity ADDSUBMAX_PL_vlg_vec_tst is
end ADDSUBMAX_PL_vlg_vec_tst;
