library verilog;
use verilog.vl_types.all;
entity AU_NONPIPELINE_vlg_vec_tst is
end AU_NONPIPELINE_vlg_vec_tst;
