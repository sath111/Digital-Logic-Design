library verilog;
use verilog.vl_types.all;
entity TEST_DP_vlg_vec_tst is
end TEST_DP_vlg_vec_tst;
