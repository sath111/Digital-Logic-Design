library verilog;
use verilog.vl_types.all;
entity SRA_SB_vlg_vec_tst is
end SRA_SB_vlg_vec_tst;
