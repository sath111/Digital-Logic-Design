library verilog;
use verilog.vl_types.all;
entity DATAPATH_PL_AU_PL_vlg_vec_tst is
end DATAPATH_PL_AU_PL_vlg_vec_tst;
