library verilog;
use verilog.vl_types.all;
entity AU_PIPELINE_vlg_vec_tst is
end AU_PIPELINE_vlg_vec_tst;
