library verilog;
use verilog.vl_types.all;
entity TEST_RISC_vlg_vec_tst is
end TEST_RISC_vlg_vec_tst;
