library verilog;
use verilog.vl_types.all;
entity PIPELINE_DP_AU_vlg_vec_tst is
end PIPELINE_DP_AU_vlg_vec_tst;
