library verilog;
use verilog.vl_types.all;
entity DATAPATH_AU_PIPELINE_vlg_vec_tst is
end DATAPATH_AU_PIPELINE_vlg_vec_tst;
