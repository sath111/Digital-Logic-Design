library verilog;
use verilog.vl_types.all;
entity CONTROLLER_vlg_vec_tst is
end CONTROLLER_vlg_vec_tst;
