library verilog;
use verilog.vl_types.all;
entity SRA_MR_vlg_vec_tst is
end SRA_MR_vlg_vec_tst;
